////////////////////////////////////////////////////////////////////////////////
// Ingress MAC Module
// Author: Niankun Rao
// Date: 2022/02/06
// Overview:
//   This module processes the incoming Ethernet byte stream, executes Layer 2
// inspection and outputs the valid Ethernet frame to the core switch fabric.
//
// Details:
//   This module executes the following Layer 2 inspections of the incoming
// Ethernet frames:
//   1. Frame statistics:
//      total octets
//      total frames (including valid and invalid frames)
//      bad CRC frames
//      under-sized frames (size < 64-byte but good CRC)
//      over-sized frames (size > MTU byte but good CRC)
//      valid frames (valid size, good CRC):
//        broadcast frames
//        multicast frames
//        unicast frames
//   2. 802.1q VLAN processing:
//      VLAN-unaware mode: all tagged and untagged frames are accepted.
//      VLAN-aware mode: Untagged frames are accepted and internally tagged with
//                       the default VLAN ID = 1.
//                       Tagged frames whose VLAN ID is in the VLAN list are
//                       accepted.
//
// Generic Table:
// +////////////////////////////////////////////////////////////////////////////
// | Generic name    | Data Type | Default Value
// |////////////////////////////////////////////////////////////////////////////
// | Description
// +////////////////////////////////////////////////////////////////////////////
//
// Port Table:
// +////////////////////////////////////////////////////////////////////////////
// | Port name       | Direction | Size, in bits | Domain      | Sense       |
// |////////////////////////////////////////////////////////////////////////////
// | Description
// +////////////////////////////////////////////////////////////////////////////
// +////////////////////////////////////////////////////////////////////////////
// | reset           | input     | 1-bit         | N/A         | active high |
// |////////////////////////////////////////////////////////////////////////////
// | Set signal to high to reset this module
// +////////////////////////////////////////////////////////////////////////////
// +////////////////////////////////////////////////////////////////////////////
// | lcl_clk         | input     | 1-bit         | N/A         | rising_edge |
// |////////////////////////////////////////////////////////////////////////////
// | Local clock running at 125MHz
// +////////////////////////////////////////////////////////////////////////////
// +////////////////////////////////////////////////////////////////////////////
// | sof_in          | input     | 1-bit         | lcl_clk     | active high |
// |////////////////////////////////////////////////////////////////////////////
// | Start of frame signal. Asserted high for 1 clock cycle before the first
// | data byte of an Ethernet frame.
// +////////////////////////////////////////////////////////////////////////////
// +////////////////////////////////////////////////////////////////////////////
// | eof_in          | input     | 1-bit         | lcl_clk     | active high |
// |////////////////////////////////////////////////////////////////////////////
// | End of frame signal. Asserted high for 1 clock cycle at the last byte of
// | an Ethernet frame.
// +////////////////////////////////////////////////////////////////////////////
// +////////////////////////////////////////////////////////////////////////////
// | valid_in        | input     | 1-bit         | lcl_clk     | active high |
// |////////////////////////////////////////////////////////////////////////////
// | Data valid signal. Asserted high for 1 clock cycle if data_out is valid.
// +////////////////////////////////////////////////////////////////////////////
// +////////////////////////////////////////////////////////////////////////////
// | data_in         | input     | 8-bit         | lcl_clk     | N/A         |
// |////////////////////////////////////////////////////////////////////////////
// | Data bus output of the stream of an Ethernet frame.
// +////////////////////////////////////////////////////////////////////////////
////////////////////////////////////////////////////////////////////////////////

`ifndef INGRESS_MAC
`define INGRESS_MAC

`default_nettype none

import ethernet_pkg::*;

module ingress_mac
(
  input wire reset   ,
  input wire lcl_clk ,

  // incoming data stream
  input wire sof_in   ,
  input wire eof_in   ,
  input wire valid_in ,
  input wire [7:0] data_in  ,

  // configurations
  input wire vlan_aware ,

  // outgoing data stream
  output logic sof_out   ,
  output logic eof_out   ,
  output logic valid_out ,
  output logic [127:0] data_out
);

endmodule

`default_nettype wire

`endif // INGRESS_MAC